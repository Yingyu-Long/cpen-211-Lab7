module regfile(
	input logic clk,
	input logic rst_n,
	input logic WE,
	input logic [1:0] selA,
	input logic [1:0] selB,
	input logic [7:0] dataW,
	output logic [7:0] dataA,
	output logic [7:0] dataB
);

             logic enable;
             logic [7:0] R0,R1,R2,R3;
             logic [1:0] rA, rB;

             assign rA = selA;
             assign rB = selB;
             assign write = WE;
				 
             always_ff @( posedge enable ) begin  // write operation
                if(write) begin
                    case (rA)
                        2'b00: begin
                            R0 <= dataW;
                        end

                        2'b01: begin
                            R1 <= dataW;
                        end

                        2'b10: begin
                            R2 <= dataW;
                        end

                        2'b11: begin
                            R3 <= dataW;
                        end
                    endcase
                end
                else if(~rst_n) begin
                    R0 <= 8'b0;
                    R1 <= 8'b0;
                    R2 <= 8'b0;
                    R3 <= 8'b0;
             end
             end

                always_comb begin  // read operation
                    case (rA)
                        2'b00: begin
                            dataA = R0;
                        end
    
                        2'b01: begin
                            dataA = R1;
                        end
    
                        2'b10: begin
                            dataA = R2;
                        end
    
                        2'b11: begin
                            dataA = R3;
                        end
                    endcase
    
                    case (rB)
                        2'b00: begin
                            dataB = R0;
                        end
    
                        2'b01: begin
                            dataB = R1;
                        end
    
                        2'b10: begin
                            dataB = R2;
                        end
    
                        2'b11: begin
                            dataB = R3;
                        end
                    endcase
                end
			
endmodule

